library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.game_types.all;


entity player is
  port
    (
      clk : in std_logic
    );
  end player;

  architecture player_arch of player is

  begin

  end player_arch;
