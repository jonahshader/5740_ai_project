library ieee;
use ieee.std_logic_1164.all;

package types is
    -- Comments for constants documentation
    -- Constants can be declared here
    
    type weight_array is array(natural range <>, natural range <>) of STD_LOGIC_VECTOR(natural range <>);
    
    -- Add other type declarations as needed
    
end package types;